d
  end

endmodule
